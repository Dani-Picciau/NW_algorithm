//Top module di tutti i blocchi presenti nella  cartella