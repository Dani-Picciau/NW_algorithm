`include "Initialization_counter.v"
`include "Insertion_Counter.v" 
`include "Match_mismatch.v"
`include "Max.v"

module Signal_manager #(
    parameter N = 128
) (

);
    
endmodule