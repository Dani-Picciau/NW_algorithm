module Index_out_B #(
    parameter N=128,
    parameter BitAddr=$clog2(N+1)
)(
    //input wire clk, rst,
    input wire en_traceB, en_read,
    input wire [BitAddr-1:0] j, j_t,
    output reg [BitAddr-1:0] index
);

    always @(en_traceB, en_read ) begin
        if(en_read) index=j;
        else if(en_traceB) index=j_t;
        else index=3'b0; // cercare un indice che non faccia danno
    end
    
endmodule